module harddrive(data_write, track, sector, clock, output_hard_drive, flag_write_hd);
  input  [31:0] data_write;
  input [6:0] track;
  input [13:0] sector;
  input flag_write_hd;
  input clock;
  output [31:0] output_hard_drive;
  integer firstClock = 0;

	// Declare the hard drive variable
	reg [31:0] HD[2:0][605:0];

	always @ (posedge clock) begin
	//load instructions
	   if (firstClock==0) begin
	 	 HD[0][0] <= 32'b01010100000000000000000100000001;//Jump to #257
	 	 HD[0][1] <= 32'b01110110101000000000000000000000;//Input to r[21]
	 	 HD[0][2] <= 32'b01101010110000000000000000000000;//Loadi #0 to r[22]
	 	 HD[0][3] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][4] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][5] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][6] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][7] <= 32'b01001100000000000000000000010011;//Branch on Zero #19
	 	 HD[0][8] <= 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
	 	 HD[0][9] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][10] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][11] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][12] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][13] <= 32'b01001100000000000000000000010000;//Branch on Zero #16
	 	 HD[0][14] <= 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
	 	 HD[0][15] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][16] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][17] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][18] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][19] <= 32'b01001100000000000000000000010111;//Branch on Zero #23
	 	 HD[0][20] <= 32'b01101010110000000000000000000011;//Loadi #3 to r[22]
	 	 HD[0][21] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][22] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][23] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][24] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][25] <= 32'b01001100000000000000000000001010;//Branch on Zero #10
	 	 HD[0][26] <= 32'b01010100000000000000001101010111;//Jump to #855
	 	 HD[0][27] <= 32'b01101010110000000000000000000000;//Loadi #0 to r[22]
	 	 HD[0][28] <= 32'b10000010110000000000000000000000;//Output r[22]
	 	 HD[0][29] <= 32'b01010100000000000000000100000001;//Jump to #257
	 	 HD[0][30] <= 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
	 	 HD[0][31] <= 32'b01101010110000000000000011000000;//Loadi #192 to r[22]
	 	 HD[0][32] <= 32'b10000110111101100000000000000000;//Loadr m[r[22]] to r[23]
	 	 HD[0][33] <= 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][34] <= 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
	 	 HD[0][35] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 HD[0][36] <= 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
	 	 HD[0][37] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[0][38] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[0][39] <= 32'b01010100000000000000000100000001;//Jump to #257
	 	 HD[0][40] <= 32'b10000010111000000000000000000000;//Output r[23]
	 	 HD[0][41] <= 32'b00000110110101100000000000000010;//ADDi r[22], #2 to r[22]
	 	 HD[0][42] <= 32'b01010100000000000000000100100000;//Jump to #288
	 	 HD[0][43] <= 32'b01110110101000000000000000000000;//Input to r[21]
	 	 HD[0][44] <= 32'b01101010110000000000000000000000;//Loadi #0 to r[22]
	 	 HD[0][45] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][46] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][47] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][48] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][49] <= 32'b01001100000000000000000000001101;//Branch on Zero #13
	 	 HD[0][50] <= 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
	 	 HD[0][51] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][52] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][53] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][54] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][55] <= 32'b01001100000000000000000000001011;//Branch on Zero #11
	 	 HD[0][56] <= 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
	 	 HD[0][57] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][58] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][59] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][60] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][61] <= 32'b01001100000000000000000000000100;//Branch on Zero #4
	 	 HD[0][62] <= 32'b01010100000000000000000101010111;//Jump to #343
	 	 HD[0][63] <= 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
	 	 HD[0][64] <= 32'b10000010110000000000000000000000;//Output r[22]
	 	 HD[0][65] <= 32'b01010100000000000000000100101011;//Jump to #299
	 	 HD[0][66] <= 32'b01010100000000000000000100000001;//Jump to #257
	 	 HD[0][67] <= 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
	 	 HD[0][68] <= 32'b01101010110000000100000000000000;//Loadi #1, #0 to r[22]
	 	 HD[0][69] <= 32'b10010110111101100000000000000000;//LoadHD m[r[22]] to r[23]
	 	 HD[0][70] <= 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][71] <= 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
	 	 HD[0][72] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 HD[0][73] <= 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
	 	 HD[0][74] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[0][75] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[0][76] <= 32'b01010100000000000000000100101011;//Jump to #299
	 	 HD[0][77] <= 32'b01101010101000000000000000000001;//Loadi #1 to r[21]
	 	 HD[0][78] <= 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][79] <= 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
	 	 HD[0][80] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 HD[0][81] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[0][82] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[0][83] <= 32'b10000010111000000000000000000000;//Output r[23]
	 	 HD[0][84] <= 32'b00000110110101100000000000100000;//ADDi r[22], #32 to r[22]
	 	 HD[0][85] <= 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
	 	 HD[0][86] <= 32'b01010100000000000000000101000101;//Jump to #325
	 	 HD[0][87] <= 32'b01101010110000000000000000000011;//Loadi #3 to r[22]
	 	 HD[0][88] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][89] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][90] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][91] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][92] <= 32'b01001100000000000000000000000000;//Branch on Zero #0
	 	 HD[0][93] <= 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
	 	 HD[0][94] <= 32'b01101010110000000000000011000000;//Loadi #192 to r[22]
	 	 HD[0][95] <= 32'b10000110111101100000000000000000;//Loadr m[r[22]] to r[23]
	 	 HD[0][96] <= 32'b01011111000000001011100000000000;//SLT if r[0] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][97] <= 32'b01011111001101110000000000000000;//SLT if r[23] < r[0], r[25] = 1 else r[25] = 0
	 	 HD[0][98] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 HD[0][99] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[0][100] <= 32'b01001100000000000000000000001001;//Branch on Zero #9
	 	 HD[0][101] <= 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][102] <= 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
	 	 HD[0][103] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 HD[0][104] <= 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
	 	 HD[0][105] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[0][106] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[0][107] <= 32'b01010100000000000000000100101011;//Jump to #299
	 	 HD[0][108] <= 32'b00000110110101100000000000000010;//ADDi r[22], #2 to r[22]
	 	 HD[0][109] <= 32'b01010100000000000000000101011111;//Jump to #351
	 	 HD[0][110] <= 32'b01101010110000000100000000000000;//Loadi #1, #0 to r[22]
	 	 HD[0][111] <= 32'b10010110111101100000000000000000;//LoadHD m[r[22]] to r[23]
	 	 HD[0][112] <= 32'b01011111000000001011100000000000;//SLT if r[0] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][113] <= 32'b01011111001101110000000000000000;//SLT if r[23] < r[0], r[25] = 1 else r[25] = 0
	 	 HD[0][114] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 HD[0][115] <= 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
	 	 HD[0][116] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[0][117] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[0][118] <= 32'b01010100000000000000000100101011;//Jump to #299
	 	 HD[0][119] <= 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][120] <= 32'b01011111001101111010100000000000;//SLT if r[23] < r[21], r[25] = 1 else r[25] = 0
	 	 HD[0][121] <= 32'b00100111001110001100100000000000;//OR r[24],r[25] to r[25]
	 	 HD[0][122] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[0][123] <= 32'b01001100000000000000000000000010;//Branch on Zero #2
	 	 HD[0][124] <= 32'b00000110110101100000000000100000;//ADDi r[22], #32 to r[22]
	 	 HD[0][125] <= 32'b01010100000000000000000101101111;//Jump to #367
	 	 HD[0][126] <= 32'b01100110101000000000000011101010;//Store r[21] in m[#234]
	 	 HD[0][127] <= 32'b01110110101000000000000000000000;//Input to r[21]
	 	 HD[0][128] <= 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
	 	 HD[0][129] <= 32'b01011110111101010000000000000000;//SLT if r[21] < r[0], r[23] = 1 else r[23] = 0
	 	 HD[0][130] <= 32'b01011111000000001010100000000000;//SLT if r[0] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][131] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][132] <= 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
	 	 HD[0][133] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][134] <= 32'b01001100000000000000000000000011;//Branch on Zero #3
	 	 HD[0][135] <= 32'b01100010110000000000000011101010;//Load m[#234] to r[22]
	 	 HD[0][136] <= 32'b10000010110000000000000000000000;//Output r[22]
	 	 HD[0][137] <= 32'b01010100000000000000000101111111;//Jump to #383
	 	 HD[0][138] <= 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
	 	 HD[0][139] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][140] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][141] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][142] <= 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
	 	 HD[0][143] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][144] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[0][145] <= 32'b01010100000000000000000100101011;//Jump to #299
	 	 HD[0][146] <= 32'b01010100000000000000001001011110;//Jump to #606
	 	 HD[0][147] <= 32'b01101011011000000000001001000110;//Loadi #582 to r[27]
	 	 HD[0][148] <= 32'b01010100000000000000000110010101;//Jump to #405
	 	 HD[0][149] <= 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
	 	 HD[0][150] <= 32'b01100100000000000000000011100000;//Store r[0] in m[#224]
	 	 HD[0][151] <= 32'b01100100000000000000000011100010;//Store r[0] in m[#226]
	 	 HD[0][152] <= 32'b01101010101000000000000011000000;//Loadi #192 to r[21]
	 	 HD[0][153] <= 32'b01100110101000000000000011100011;//Store r[21] in m[#227]
	 	 HD[0][154] <= 32'b01100010101000000000000011100011;//Load m[#227] to r[21]
	 	 HD[0][155] <= 32'b10000110110101010000000000000000;//Loadr m[r[21]] to r[22]
	 	 HD[0][156] <= 32'b01011110111101100000000000000000;//SLT if r[22] < r[0], r[23] = 1 else r[23] = 0
	 	 HD[0][157] <= 32'b01011111000000001011000000000000;//SLT if r[0] < r[22], r[24] = 1 else r[24] = 0
	 	 HD[0][158] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][159] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][160] <= 32'b01001100000000000000000000010100;//Branch on Zero #20
	 	 HD[0][161] <= 32'b01101011000000000000000000000001;//Loadi #1 to r[24]
	 	 HD[0][162] <= 32'b01011111000110001011000000000000;//SLT if r[24] < r[22], r[24] = 1 else r[24] = 0
	 	 HD[0][163] <= 32'b01111100000110000000000000000000;//Pre Branch r[24]
	 	 HD[0][164] <= 32'b01001100000000000000000000001100;//Branch on Zero #12
	 	 HD[0][165] <= 32'b01100010101000000000000011100011;//Load m[#227] to r[21]
	 	 HD[0][166] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][167] <= 32'b10000110110101010000000000000000;//Loadr m[r[21]] to r[22]
	 	 HD[0][168] <= 32'b01011110111101100000000000000000;//SLT if r[22] < r[0], r[23] = 1 else r[23] = 0
	 	 HD[0][169] <= 32'b01011111000000001011000000000000;//SLT if r[0] < r[22], r[24] = 1 else r[24] = 0
	 	 HD[0][170] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][171] <= 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
	 	 HD[0][172] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][173] <= 32'b01001100000000000000000000000011;//Branch on Zero #3
	 	 HD[0][174] <= 32'b01100011000000000000000011100010;//Load m[#226] to r[24]
	 	 HD[0][175] <= 32'b00000111000110000000000000000001;//ADDi r[24], #1 to r[24]
	 	 HD[0][176] <= 32'b01100111000000000000000011100010;//Store r[24] in m[#226]
	 	 HD[0][177] <= 32'b01100010101000000000000011100011;//Load m[#227] to r[21]
	 	 HD[0][178] <= 32'b00000110101101010000000000000010;//ADDi r[21], #2 to r[21]
	 	 HD[0][179] <= 32'b01100110101000000000000011100011;//Store r[21] in m[#227]
	 	 HD[0][180] <= 32'b01010100000000000000000110011010;//Jump to #410
	 	 HD[0][181] <= 32'b01100010101000000000000011100010;//Load m[#226] to r[21]
	 	 HD[0][182] <= 32'b01101010110000000000000000000010;//Loadi #2 to r[22]
	 	 HD[0][183] <= 32'b01011110110101101010100000000000;//SLT if r[22] < r[21], r[22] = 1 else r[22] = 0
	 	 HD[0][184] <= 32'b01111100000101100000000000000000;//Pre Branch r[22]
	 	 HD[0][185] <= 32'b01001100000000000000000000000010;//Branch on Zero #2
	 	 HD[0][186] <= 32'b01101010101000000000000000000001;//Loadi #1 to r[21]
	 	 HD[0][187] <= 32'b01100110101000000000000011100000;//Store r[21] in m[#224]
	 	 HD[0][188] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][189] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][190] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][191] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][192] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][193] <= 32'b10001100000110110000000000000000;//Jump to r[27]
	 	 HD[0][194] <= 32'b01100010101000000000000001100000;//Load m[#96] to r[21]
	 	 HD[0][195] <= 32'b10000010101000000000000000000000;//Output r[21]
	 	 HD[0][196] <= 32'b01101011011000000000000111110000;//Loadi #496 to r[27]
	 	 HD[0][197] <= 32'b01100010101000000000000011101010;//Load m[#234] to r[21]
	 	 HD[0][198] <= 32'b01100110101000000000000011100100;//Store r[21] in m[#228]
	 	 HD[0][199] <= 32'b01100100000000000000000011100101;//Store r[0] in m[#229]
	 	 HD[0][200] <= 32'b01100100000000000000000011100110;//Store r[0] in m[#230]
	 	 HD[0][201] <= 32'b01101010101000000000000000000001;//Loadi #1 to r[21]
	 	 HD[0][202] <= 32'b01100110101000000000000011100111;//Store r[21] in m[#231]
	 	 HD[0][203] <= 32'b01100100000000000000000011101000;//Store r[0] in m[#232]
	 	 HD[0][204] <= 32'b01010100000000000000000111001101;//Jump to #461
	 	 HD[0][205] <= 32'b01101010101000000100000000000000;//Loadi #1, #0 to r[21]
	 	 HD[0][206] <= 32'b01100110101000000000000011101001;//Store r[21] in m[#233]
	 	 HD[0][207] <= 32'b01100010101000000000000011101001;//Load m[#233] to r[21]
	 	 HD[0][208] <= 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
	 	 HD[0][209] <= 32'b01100010111000000000000011100100;//Load m[#228] to r[23]
	 	 HD[0][210] <= 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][211] <= 32'b01011111001101111011000000000000;//SLT if r[23] < r[22], r[25] = 1 else r[25] = 0
	 	 HD[0][212] <= 32'b00100111000110001100100000000000;//OR r[24],r[25] to r[24]
	 	 HD[0][213] <= 32'b01111100000110000000000000000000;//Pre Branch r[24]
	 	 HD[0][214] <= 32'b01001100000000000000000000000010;//Branch on Zero #2
	 	 HD[0][215] <= 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
	 	 HD[0][216] <= 32'b01010100000000000000000111001110;//Jump to #462
	 	 HD[0][217] <= 32'b01100010101000000000000011101001;//Load m[#233] to r[21]
	 	 HD[0][218] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][219] <= 32'b01100010110000000000000011100101;//Load m[#229] to r[22]
	 	 HD[0][220] <= 32'b10010010110101010000000000000000;//hdStore r[22] in m[r[21]] 
	 	 HD[0][221] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][222] <= 32'b01100010110000000000000011100110;//Load m[#230] to r[22]
	 	 HD[0][223] <= 32'b10010010110101010000000000000000;//hdStore r[22] in m[r[21]] 
	 	 HD[0][224] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][225] <= 32'b01100010110000000000000011100111;//Load m[#231] to r[22]
	 	 HD[0][226] <= 32'b10010010110101010000000000000000;//hdStore r[22] in m[r[21]] 
	 	 HD[0][227] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][228] <= 32'b01100010110000000000000011101000;//Load m[#232] to r[22]
	 	 HD[0][229] <= 32'b10010010110101010000000000000000;//hdStore r[22] in m[r[21]] 
	 	 HD[0][230] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][231] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][232] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][233] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][234] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][235] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][236] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][237] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][238] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][239] <= 32'b10001100000110110000000000000000;//Jump to r[27]
	 	 HD[0][240] <= 32'b01101011011000000000001000001110;//Loadi #526 to r[27]
	 	 HD[0][241] <= 32'b01100010101000000000000011101010;//Load m[#234] to r[21]
	 	 HD[0][242] <= 32'b01100110101000000000000011101011;//Store r[21] in m[#235]
	 	 HD[0][243] <= 32'b01100100000000000000000011101100;//Store r[0] in m[#236]
	 	 HD[0][244] <= 32'b01010100000000000000000111110101;//Jump to #501
	 	 HD[0][245] <= 32'b01101010101000000000000011000000;//Loadi #192 to r[21]
	 	 HD[0][246] <= 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
	 	 HD[0][247] <= 32'b10000111000101010000000000000000;//Loadr m[r[21]] to r[24]
	 	 HD[0][248] <= 32'b01011110111101101100000000000000;//SLT if r[22] < r[24], r[23] = 1 else r[23] = 0
	 	 HD[0][249] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][250] <= 32'b01001100000000000000000000000010;//Branch on Zero #2
	 	 HD[0][251] <= 32'b00000110101101010000000000000010;//ADDi r[21], #2 to r[21]
	 	 HD[0][252] <= 32'b01010100000000000000000111110111;//Jump to #503
	 	 HD[0][253] <= 32'b01100010110000000000000011101011;//Load m[#235] to r[22]
	 	 HD[0][254] <= 32'b01100010111000000000000011101100;//Load m[#236] to r[23]
	 	 HD[0][255] <= 32'b10001010110101010000000000000000;//rStore r[22] in m[r[21]] 
	 	 HD[0][256] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][257] <= 32'b10001010111101010000000000000000;//rStore r[23] in m[r[21]] 
	 	 HD[0][258] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][259] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][260] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][261] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][262] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][263] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][264] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][265] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][266] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][267] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][268] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][269] <= 32'b10001100000110110000000000000000;//Jump to r[27]
	 	 HD[0][270] <= 32'b01100010101000000000000011101010;//Load m[#234] to r[21]
	 	 HD[0][271] <= 32'b01100110101000000000000011110001;//Store r[21] in m[#241]
	 	 HD[0][272] <= 32'b01101011011000000000001000101011;//Loadi #555 to r[27]
	 	 HD[0][273] <= 32'b10000010101000000000000000000000;//Output r[21]
	 	 HD[0][274] <= 32'b01101010110000000100000000000000;//Loadi #1, #0 to r[22]
	 	 HD[0][275] <= 32'b01100110110000000000000011110011;//Store r[22] in m[#243]
	 	 HD[0][276] <= 32'b01100010101000000000000011110011;//Load m[#243] to r[21]
	 	 HD[0][277] <= 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
	 	 HD[0][278] <= 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][279] <= 32'b01011111000101100000000000000000;//SLT if r[22] < r[0], r[24] = 1 else r[24] = 0
	 	 HD[0][280] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][281] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][282] <= 32'b01001100000000000000000000001110;//Branch on Zero #14
	 	 HD[0][283] <= 32'b01100011001000000000000011110001;//Load m[#241] to r[25]
	 	 HD[0][284] <= 32'b01011110111101101100100000000000;//SLT if r[22] < r[25], r[23] = 1 else r[23] = 0
	 	 HD[0][285] <= 32'b01011111000110011011000000000000;//SLT if r[25] < r[22], r[24] = 1 else r[24] = 0
	 	 HD[0][286] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][287] <= 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
	 	 HD[0][288] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][289] <= 32'b01001100000000000000000000000100;//Branch on Zero #4
	 	 HD[0][290] <= 32'b00000110110101010000000000000101;//ADDi r[21], #5 to r[22]
	 	 HD[0][291] <= 32'b10010110110101100000000000000000;//LoadHD m[r[22]] to r[22]
	 	 HD[0][292] <= 32'b01100110110000000000000011110010;//Store r[22] in m[#242]
	 	 HD[0][293] <= 32'b01010100000000000000001000101010;//Jump to #554
	 	 HD[0][294] <= 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
	 	 HD[0][295] <= 32'b01100110101000000000000011110011;//Store r[21] in m[#243]
	 	 HD[0][296] <= 32'b01010100000000000000001000010100;//Jump to #532
	 	 HD[0][297] <= 32'b01100100000000000000000011110010;//Store r[0] in m[#242]
	 	 HD[0][298] <= 32'b10001100000110110000000000000000;//Jump to r[27]
	 	 HD[0][299] <= 32'b01100010101000000000000011110010;//Load m[#242] to r[21]
	 	 HD[0][300] <= 32'b01100110101000000000000011101110;//Store r[21] in m[#238]
	 	 HD[0][301] <= 32'b01101011011000000000001001000101;//Loadi #581 to r[27]
	 	 HD[0][302] <= 32'b01100100000000000000000011101111;//Store r[0] in m[#239]
	 	 HD[0][303] <= 32'b01101010101000000000000001000000;//Loadi #64 to r[21]
	 	 HD[0][304] <= 32'b01100010110000000000000011101110;//Load m[#238] to r[22]
	 	 HD[0][305] <= 32'b00010010101101011011000000000000;//TIMES r[21],r[22] to r[21]
	 	 HD[0][306] <= 32'b10000010110000000000000000000000;//Output r[22]
	 	 HD[0][307] <= 32'b01101010110000001000000000000000;//Loadi #2, #0 to r[22]
	 	 HD[0][308] <= 32'b00000010101101011011000000000000;//ADD r[21],r[22] to r[21]
	 	 HD[0][309] <= 32'b01100110101000000000000011110000;//Store r[21] in m[#240]
	 	 HD[0][310] <= 32'b01100010101000000000000011110000;//Load m[#240] to r[21]
	 	 HD[0][311] <= 32'b01100010110000000000000011101111;//Load m[#239] to r[22]
	 	 HD[0][312] <= 32'b00000010101101011011000000000000;//ADD r[21],r[22] to r[21]
	 	 HD[0][313] <= 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
	 	 HD[0][314] <= 32'b01011110111101100000000000000000;//SLT if r[22] < r[0], r[23] = 1 else r[23] = 0
	 	 HD[0][315] <= 32'b01011111000000001011000000000000;//SLT if r[0] < r[22], r[24] = 1 else r[24] = 0
	 	 HD[0][316] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][317] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][318] <= 32'b01001100000000000000000000000101;//Branch on Zero #5
	 	 HD[0][319] <= 32'b01100010111000000000000011101111;//Load m[#239] to r[23]
	 	 HD[0][320] <= 32'b10011010110101110000000000000000;//rStore r[22] in m[r[23]] 
	 	 HD[0][321] <= 32'b00000110111101110000000000000001;//ADDi r[23], #1 to r[23]
	 	 HD[0][322] <= 32'b01100110111000000000000011101111;//Store r[23] in m[#239]
	 	 HD[0][323] <= 32'b01010100000000000000001000110110;//Jump to #566
	 	 HD[0][324] <= 32'b10001100000110110000000000000000;//Jump to r[27]
	 	 HD[0][325] <= 32'b01010100000000000000000000000000;//Jump to #0
	 	 HD[0][326] <= 32'b01101011011000000000001001010110;//Loadi #598 to r[27]
	 	 HD[0][327] <= 32'b01010100000000000000001001001000;//Jump to #584
	 	 HD[0][328] <= 32'b01100100000000000000000011110100;//Store r[0] in m[#244]
	 	 HD[0][329] <= 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
	 	 HD[0][330] <= 32'b01101010101000000000000011000000;//Loadi #192 to r[21]
	 	 HD[0][331] <= 32'b10000110111101010000000000000000;//Loadr m[r[21]] to r[23]
	 	 HD[0][332] <= 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][333] <= 32'b01111100000110000000000000000000;//Pre Branch r[24]
	 	 HD[0][334] <= 32'b01001100000000000000000000000100;//Branch on Zero #4
	 	 HD[0][335] <= 32'b01101011001000000000000000000001;//Loadi #1 to r[25]
	 	 HD[0][336] <= 32'b01100111001000000000000011110100;//Store r[25] in m[#244]
	 	 HD[0][337] <= 32'b00000110101101010000000000000010;//ADDi r[21], #2 to r[21]
	 	 HD[0][338] <= 32'b01010100000000000000001001001011;//Jump to #587
	 	 HD[0][339] <= 32'b01101010100000000000000111000010;//Loadi #450 to r[20]
	 	 HD[0][340] <= 32'b10000010100000000000000000000000;//Output r[20]
	 	 HD[0][341] <= 32'b10001100000110110000000000000000;//Jump to r[27]
	 	 HD[0][342] <= 32'b01100010101000000000000011110100;//Load m[#244] to r[21]
	 	 HD[0][343] <= 32'b01011110110101010000000000000000;//SLT if r[21] < r[0], r[22] = 1 else r[22] = 0
	 	 HD[0][344] <= 32'b01011110111000001010100000000000;//SLT if r[0] < r[21], r[23] = 1 else r[23] = 0
	 	 HD[0][345] <= 32'b00100110110101101011100000000000;//OR r[22],r[23] to r[22]
	 	 HD[0][346] <= 32'b00110110110101100000000000000000;//NOT r[22] to r[22]
	 	 HD[0][347] <= 32'b01111100000101100000000000000000;//Pre Branch r[22]
	 	 HD[0][348] <= 32'b01001100000000000000000000011011;//Branch on Zero #27
	 	 HD[0][349] <= 32'b01010100000000000000000111000100;//Jump to #452
	 	 HD[0][350] <= 32'b01101010110000000000000000000001;//Loadi #1 to r[22]
	 	 HD[0][351] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][352] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][353] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][354] <= 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
	 	 HD[0][355] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][356] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[0][357] <= 32'b01010100000000000000001001000110;//Jump to #582
	 	 HD[0][358] <= 32'b01101010110000000000000000000011;//Loadi #3 to r[22]
	 	 HD[0][359] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][360] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][361] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][362] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][363] <= 32'b01001100000000000000000000000000;//Branch on Zero #0
	 	 HD[0][364] <= 32'b01101010110000000000000000000100;//Loadi #4 to r[22]
	 	 HD[0][365] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][366] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][367] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][368] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][369] <= 32'b01001100000000000000000000000000;//Branch on Zero #0
	 	 HD[0][370] <= 32'b01101010110000000000000000000101;//Loadi #5 to r[22]
	 	 HD[0][371] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][372] <= 32'b01011111000101101010100000000000;//SLT if r[22] < r[21], r[24] = 1 else r[24] = 0
	 	 HD[0][373] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][374] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][375] <= 32'b01001100000000000000000000000000;//Branch on Zero #0
	 	 HD[0][376] <= 32'b01101011011000000000001001111010;//Loadi #634 to r[27]
	 	 HD[0][377] <= 32'b01101010100000000000000111000011;//Loadi #451 to r[20]
	 	 HD[0][378] <= 32'b10000010100000000000000000000000;//Output r[20]
	 	 HD[0][379] <= 32'b01101010100000000000000111000100;//Loadi #452 to r[20]
	 	 HD[0][380] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][381] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][382] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][383] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][384] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][385] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[0][386] <= 32'b01101011011000000000001010100110;//Loadi #678 to r[27]
	 	 HD[0][387] <= 32'b01101010101000000100000000000000;//Loadi #1, #0 to r[21]
	 	 HD[0][388] <= 32'b01100110101000000000000011110110;//Store r[21] in m[#246]
	 	 HD[0][389] <= 32'b01100010101000000000000011110110;//Load m[#246] to r[21]
	 	 HD[0][390] <= 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
	 	 HD[0][391] <= 32'b01011110111101100000000000000000;//SLT if r[22] < r[0], r[23] = 1 else r[23] = 0
	 	 HD[0][392] <= 32'b01011111000000001011000000000000;//SLT if r[0] < r[22], r[24] = 1 else r[24] = 0
	 	 HD[0][393] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][394] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][395] <= 32'b01001100000000000000000000011001;//Branch on Zero #25
	 	 HD[0][396] <= 32'b01101011000000000000000000000001;//Loadi #1 to r[24]
	 	 HD[0][397] <= 32'b01011111001101101100000000000000;//SLT if r[22] < r[24], r[25] = 1 else r[25] = 0
	 	 HD[0][398] <= 32'b01011111000110001011000000000000;//SLT if r[24] < r[22], r[24] = 1 else r[24] = 0
	 	 HD[0][399] <= 32'b00100111000110001100100000000000;//OR r[24],r[25] to r[24]
	 	 HD[0][400] <= 32'b01111100000110000000000000000000;//Pre Branch r[24]
	 	 HD[0][401] <= 32'b01001100000000000000000000010000;//Branch on Zero #16
	 	 HD[0][402] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][403] <= 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
	 	 HD[0][404] <= 32'b01011111001000001011100000000000;//SLT if r[0] < r[23], r[25] = 1 else r[25] = 0
	 	 HD[0][405] <= 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
	 	 HD[0][406] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[0][407] <= 32'b01001100000000000000000000001010;//Branch on Zero #10
	 	 HD[0][408] <= 32'b00000110101101010000000000000010;//ADDi r[21], #2 to r[21]
	 	 HD[0][409] <= 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
	 	 HD[0][410] <= 32'b01101011000000000000000000000001;//Loadi #1 to r[24]
	 	 HD[0][411] <= 32'b01011111001110001011100000000000;//SLT if r[24] < r[23], r[25] = 1 else r[25] = 0
	 	 HD[0][412] <= 32'b01011111010101111100000000000000;//SLT if r[23] < r[24], r[26] = 1 else r[26] = 0
	 	 HD[0][413] <= 32'b00100111001110011101000000000000;//OR r[25],r[26] to r[25]
	 	 HD[0][414] <= 32'b00110111001110010000000000000000;//NOT r[25] to r[25]
	 	 HD[0][415] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[0][416] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[0][417] <= 32'b01100110110000000000000011110111;//Store r[22] in m[#247]
	 	 HD[0][418] <= 32'b01100010101000000000000011110110;//Load m[#246] to r[21]
	 	 HD[0][419] <= 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
	 	 HD[0][420] <= 32'b01010100000000000000001010000100;//Jump to #644
	 	 HD[0][421] <= 32'b10001100000110110000000000000000;//Jump to r[27]
	 	 HD[0][422] <= 32'b01101011011000000000001011100001;//Loadi #737 to r[27]
	 	 HD[0][423] <= 32'b10000010100000000000000000000000;//Output r[20]
	 	 HD[0][424] <= 32'b01101010101000000000000010100000;//Loadi #160 to r[21]
	 	 HD[0][425] <= 32'b01101010110000000000000010101010;//Loadi #170 to r[22]
	 	 HD[0][426] <= 32'b01100110101000000000000011111000;//Store r[21] in m[#248]
	 	 HD[0][427] <= 32'b01100010101000000000000011111000;//Load m[#248] to r[21]
	 	 HD[0][428] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][429] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][430] <= 32'b01001100000000000000000000000011;//Branch on Zero #3
	 	 HD[0][431] <= 32'b10001000000101010000000000000000;//rStore r[0] in m[r[21]] 
	 	 HD[0][432] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][433] <= 32'b01010100000000000000001010101010;//Jump to #682
	 	 HD[0][434] <= 32'b01101010101000000100000000000000;//Loadi #1, #0 to r[21]
	 	 HD[0][435] <= 32'b01100110101000000000000011111000;//Store r[21] in m[#248]
	 	 HD[0][436] <= 32'b01100010101000000000000011111000;//Load m[#248] to r[21]
	 	 HD[0][437] <= 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
	 	 HD[0][438] <= 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][439] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][440] <= 32'b01001100000000000000000000010110;//Branch on Zero #22
	 	 HD[0][441] <= 32'b01101011000000000000000000000001;//Loadi #1 to r[24]
	 	 HD[0][442] <= 32'b01011110111101101100000000000000;//SLT if r[22] < r[24], r[23] = 1 else r[23] = 0
	 	 HD[0][443] <= 32'b01011111001110001011000000000000;//SLT if r[24] < r[22], r[25] = 1 else r[25] = 0
	 	 HD[0][444] <= 32'b00100110111101111100100000000000;//OR r[23],r[25] to r[23]
	 	 HD[0][445] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][446] <= 32'b01001100000000000000000000001101;//Branch on Zero #13
	 	 HD[0][447] <= 32'b00000110101101010000000000000011;//ADDi r[21], #3 to r[21]
	 	 HD[0][448] <= 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
	 	 HD[0][449] <= 32'b01011110111101101100000000000000;//SLT if r[22] < r[24], r[23] = 1 else r[23] = 0
	 	 HD[0][450] <= 32'b01011111001110001011000000000000;//SLT if r[24] < r[22], r[25] = 1 else r[25] = 0
	 	 HD[0][451] <= 32'b00100110111101111100100000000000;//OR r[23],r[25] to r[23]
	 	 HD[0][452] <= 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
	 	 HD[0][453] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][454] <= 32'b01001100000000000000000000000101;//Branch on Zero #5
	 	 HD[0][455] <= 32'b01100010101000000000000011111000;//Load m[#248] to r[21]
	 	 HD[0][456] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][457] <= 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
	 	 HD[0][458] <= 32'b00000110110101100000000010100000;//ADDi r[22], #160 to r[22]
	 	 HD[0][459] <= 32'b10001011000101100000000000000000;//rStore r[24] in m[r[22]] 
	 	 HD[0][460] <= 32'b01100010101000000000000011111000;//Load m[#248] to r[21]
	 	 HD[0][461] <= 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
	 	 HD[0][462] <= 32'b01010100000000000000001010110011;//Jump to #691
	 	 HD[0][463] <= 32'b01101010101000000000000010100000;//Loadi #160 to r[21]
	 	 HD[0][464] <= 32'b01101010110000000000000010101010;//Loadi #170 to r[22]
	 	 HD[0][465] <= 32'b01100110101000000000000011111000;//Store r[21] in m[#248]
	 	 HD[0][466] <= 32'b01100010101000000000000011111000;//Load m[#248] to r[21]
	 	 HD[0][467] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][468] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][469] <= 32'b01001100000000000000000000001010;//Branch on Zero #10
	 	 HD[0][470] <= 32'b10000110111101010000000000000000;//Loadr m[r[21]] to r[23]
	 	 HD[0][471] <= 32'b01011110111000001011100000000000;//SLT if r[0] < r[23], r[23] = 1 else r[23] = 0
	 	 HD[0][472] <= 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
	 	 HD[0][473] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][474] <= 32'b01001100000000000000000000000011;//Branch on Zero #3
	 	 HD[0][475] <= 32'b00001110101101010000000010100000;//SUBi r[21], #160 to r[21]
	 	 HD[0][476] <= 32'b01100110101000000000000011111001;//Store r[21] in m[#249]
	 	 HD[0][477] <= 32'b01010100000000000000001011100000;//Jump to #736
	 	 HD[0][478] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][479] <= 32'b01010100000000000000001011010001;//Jump to #721
	 	 HD[0][480] <= 32'b10001100000110110000000000000000;//Jump to r[27]
	 	 HD[0][481] <= 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
	 	 HD[0][482] <= 32'b01100110101000000000000011111010;//Store r[21] in m[#250]
	 	 HD[0][483] <= 32'b01100010101000000000000011111001;//Load m[#249] to r[21]
	 	 HD[0][484] <= 32'b01100110101000000000000011111011;//Store r[21] in m[#251]
	 	 HD[0][485] <= 32'b01101011011000000000001100010100;//Loadi #788 to r[27]
	 	 HD[0][486] <= 32'b10000010100000000000000000000000;//Output r[20]
	 	 HD[0][487] <= 32'b01101010101000000100000000000000;//Loadi #1, #0 to r[21]
	 	 HD[0][488] <= 32'b01100110101000000000000011111100;//Store r[21] in m[#252]
	 	 HD[0][489] <= 32'b01100010101000000000000011111100;//Load m[#252] to r[21]
	 	 HD[0][490] <= 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
	 	 HD[0][491] <= 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][492] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][493] <= 32'b01001100000000000000000000010000;//Branch on Zero #16
	 	 HD[0][494] <= 32'b01100010111000000000000011111010;//Load m[#250] to r[23]
	 	 HD[0][495] <= 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][496] <= 32'b01011110111101111011000000000000;//SLT if r[23] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][497] <= 32'b00100110111101111100000000000000;//OR r[23],r[24] to r[23]
	 	 HD[0][498] <= 32'b00110110111101110000000000000000;//NOT r[23] to r[23]
	 	 HD[0][499] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][500] <= 32'b01001100000000000000000000000110;//Branch on Zero #6
	 	 HD[0][501] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][502] <= 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
	 	 HD[0][503] <= 32'b01100110111000000000000011111101;//Store r[23] in m[#253]
	 	 HD[0][504] <= 32'b01100010111000000000000011111011;//Load m[#251] to r[23]
	 	 HD[0][505] <= 32'b10010010111101010000000000000000;//hdStore r[23] in m[r[21]] 
	 	 HD[0][506] <= 32'b01010100000000000000001011111110;//Jump to #766
	 	 HD[0][507] <= 32'b01100010101000000000000011111100;//Load m[#252] to r[21]
	 	 HD[0][508] <= 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
	 	 HD[0][509] <= 32'b01010100000000000000001011101000;//Jump to #744
	 	 HD[0][510] <= 32'b01100010110000000000000011111101;//Load m[#253] to r[22]
	 	 HD[0][511] <= 32'b01101010111000000000000001000000;//Loadi #64 to r[23]
	 	 HD[0][512] <= 32'b00010010110101101011100000000000;//TIMES r[22],r[23] to r[22]
	 	 HD[0][513] <= 32'b01100110110000000000000011111101;//Store r[22] in m[#253]
	 	 HD[0][514] <= 32'b01100010110000000000000011111011;//Load m[#251] to r[22]
	 	 HD[0][515] <= 32'b00010010110101101011100000000000;//TIMES r[22],r[23] to r[22]
	 	 HD[0][516] <= 32'b01100110110000000000000011111110;//Store r[22] in m[#254]
	 	 HD[0][517] <= 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
	 	 HD[0][518] <= 32'b01100110101000000000000011111100;//Store r[21] in m[#252]
	 	 HD[0][519] <= 32'b01100010101000000000000011111100;//Load m[#252] to r[21]
	 	 HD[0][520] <= 32'b01011111000101011011100000000000;//SLT if r[21] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][521] <= 32'b01111100000110000000000000000000;//Pre Branch r[24]
	 	 HD[0][522] <= 32'b01001100000000000000000000001000;//Branch on Zero #8
	 	 HD[0][523] <= 32'b01100010110000000000000011111101;//Load m[#253] to r[22]
	 	 HD[0][524] <= 32'b00000010110101011011000000000000;//ADD r[21],r[22] to r[22]
	 	 HD[0][525] <= 32'b10000110110101100000000000000000;//Loadr m[r[22]] to r[22]
	 	 HD[0][526] <= 32'b01100011000000000000000011111110;//Load m[#254] to r[24]
	 	 HD[0][527] <= 32'b00000011000101011100000000000000;//ADD r[21],r[24] to r[24]
	 	 HD[0][528] <= 32'b10001010110110000000000000000000;//rStore r[22] in m[r[24]] 
	 	 HD[0][529] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][530] <= 32'b01010100000000000000001100000110;//Jump to #774
	 	 HD[0][531] <= 32'b10001100000110110000000000000000;//Jump to r[27]
	 	 HD[0][532] <= 32'b01100010101000000000000011110111;//Load m[#247] to r[21]
	 	 HD[0][533] <= 32'b01100110101000000000000011111111;//Store r[21] in m[#255]
	 	 HD[0][534] <= 32'b01101011011000000000000111000100;//Loadi #452 to r[27]
	 	 HD[0][535] <= 32'b10000010100000000000000000000000;//Output r[20]
	 	 HD[0][536] <= 32'b01101010101000000100000000000000;//Loadi #1, #0 to r[21]
	 	 HD[0][537] <= 32'b01100110101000000000000100000000;//Store r[21] in m[#256]
	 	 HD[0][538] <= 32'b01100010101000000000000100000000;//Load m[#256] to r[21]
	 	 HD[0][539] <= 32'b10010110110101010000000000000000;//LoadHD m[r[21]] to r[22]
	 	 HD[0][540] <= 32'b01011110111000001011000000000000;//SLT if r[0] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[0][541] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[0][542] <= 32'b01001100000000000000000000001011;//Branch on Zero #11
	 	 HD[0][543] <= 32'b01100010111000000000000011111111;//Load m[#255] to r[23]
	 	 HD[0][544] <= 32'b01011111000101101011100000000000;//SLT if r[22] < r[23], r[24] = 1 else r[24] = 0
	 	 HD[0][545] <= 32'b01011111001101111011000000000000;//SLT if r[23] < r[22], r[25] = 1 else r[25] = 0
	 	 HD[0][546] <= 32'b00100111000110001100100000000000;//OR r[24],r[25] to r[24]
	 	 HD[0][547] <= 32'b00110111000110000000000000000000;//NOT r[24] to r[24]
	 	 HD[0][548] <= 32'b01111100000110000000000000000000;//Pre Branch r[24]
	 	 HD[0][549] <= 32'b01001100000000000000000000000001;//Branch on Zero #1
	 	 HD[0][550] <= 32'b01010100000000000000001100101010;//Jump to #810
	 	 HD[0][551] <= 32'b01100010101000000000000100000000;//Load m[#256] to r[21]
	 	 HD[0][552] <= 32'b00000110101101010000000000100000;//ADDi r[21], #32 to r[21]
	 	 HD[0][553] <= 32'b01010100000000000000001100011001;//Jump to #793
	 	 HD[0][554] <= 32'b01100110101000000000000100000000;//Store r[21] in m[#256]
	 	 HD[0][555] <= 32'b01100010101000000000000100000000;//Load m[#256] to r[21]
	 	 HD[0][556] <= 32'b00000110101101010000000000000100;//ADDi r[21], #4 to r[21]
	 	 HD[0][557] <= 32'b10010011100101010000000000000000;//hdStore r[28] in m[r[21]] 
	 	 HD[0][558] <= 32'b00000110101101010000000000001000;//ADDi r[21], #8 to r[21]
	 	 HD[0][559] <= 32'b10010000000101010000000000000000;//hdStore r[0] in m[r[21]] 
	 	 HD[0][560] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][561] <= 32'b10010000001101010000000000000000;//hdStore r[1] in m[r[21]] 
	 	 HD[0][562] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][563] <= 32'b10010000010101010000000000000000;//hdStore r[2] in m[r[21]] 
	 	 HD[0][564] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][565] <= 32'b10010000011101010000000000000000;//hdStore r[3] in m[r[21]] 
	 	 HD[0][566] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][567] <= 32'b10010000100101010000000000000000;//hdStore r[4] in m[r[21]] 
	 	 HD[0][568] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][569] <= 32'b10010000101101010000000000000000;//hdStore r[5] in m[r[21]] 
	 	 HD[0][570] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][571] <= 32'b10010000110101010000000000000000;//hdStore r[6] in m[r[21]] 
	 	 HD[0][572] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][573] <= 32'b10010000111101010000000000000000;//hdStore r[7] in m[r[21]] 
	 	 HD[0][574] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][575] <= 32'b10010001000101010000000000000000;//hdStore r[8] in m[r[21]] 
	 	 HD[0][576] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][577] <= 32'b10010001001101010000000000000000;//hdStore r[9] in m[r[21]] 
	 	 HD[0][578] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][579] <= 32'b10010001010101010000000000000000;//hdStore r[10] in m[r[21]] 
	 	 HD[0][580] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][581] <= 32'b10010001011101010000000000000000;//hdStore r[11] in m[r[21]] 
	 	 HD[0][582] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][583] <= 32'b10010001100101010000000000000000;//hdStore r[12] in m[r[21]] 
	 	 HD[0][584] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][585] <= 32'b10010001101101010000000000000000;//hdStore r[13] in m[r[21]] 
	 	 HD[0][586] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][587] <= 32'b10010001110101010000000000000000;//hdStore r[14] in m[r[21]] 
	 	 HD[0][588] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][589] <= 32'b10010001111101010000000000000000;//hdStore r[15] in m[r[21]] 
	 	 HD[0][590] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][591] <= 32'b10010010000101010000000000000000;//hdStore r[16] in m[r[21]] 
	 	 HD[0][592] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][593] <= 32'b10010010001101010000000000000000;//hdStore r[17] in m[r[21]] 
	 	 HD[0][594] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][595] <= 32'b10010010010101010000000000000000;//hdStore r[18] in m[r[21]] 
	 	 HD[0][596] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[0][597] <= 32'b10010010011101010000000000000000;//hdStore r[19] in m[r[21]] 
	 	 HD[0][598] <= 32'b10001100000110110000000000000000;//Jump to r[27]
		 HD[0][599] <= 32'b00000000000000000000000000000000;
HD[1][0] <= 32'b00000000000000000000000000000001;
HD[1][32] <= 32'b00000000000000000000000000000110;
HD[1][33] <= 32'b00000000000000000000000000000111;
HD[1][34] <= 32'b00000000000000000000000000000111;
HD[1][35] <= 32'b00000000000000000000000000000111;
HD[1][37] <= 32'b00000000000000000000000000000010;
HD[1][38] <= 32'b00000000000000000000000000000111;
HD[1][64] <= 32'b00000000000000000000000000001001;
HD[1][69] <= 32'b00000000000000000000000000000000;
HD[1][96] <= 32'b00000000000000000000000000001010;
HD[1][101] <= 32'b00000000000000000000000000000001;
HD[1][128] <= 32'b00000000000000000000000000000000;
HD[2][0] <= 32'b01101100000000000000000000000000;//Nop
HD[2][1] <= 32'b01110100100000000000000000000000;//Input to r[4]
HD[2][2] <= 32'b01110100101000000000000000000000;//Input to r[5]
HD[2][3] <= 32'b01100100100000000000000000001000;//Store r[4] in m[#8]
HD[2][4] <= 32'b01100000110000000000000000001000;//Load m[#8] to r[6]
HD[2][5] <= 32'b00000000111001000010100000000000;//ADD r[4],r[5] to r[7]
HD[2][6] <= 32'b10000000111000000000000000000000;//Output r[7]
HD[2][7] <= 32'b01110000000000000000000000000000;//Hlt
HD[2][8] <= 32'b00000000000000000000000000000000;
HD[2][64] <= 32'b01101100000000000000000000000000;//Nop
HD[2][65] <= 32'b01110100100000000000000000000000;//Input to r[4]
HD[2][66] <= 32'b01110100101000000000000000000000;//Input to r[5]
HD[2][67] <= 32'b01100100100000000000000000001000;//Store r[4] in m[#8]
HD[2][68] <= 32'b01100000110000000000000000001000;//Load m[#8] to r[6]
HD[2][69] <= 32'b00001000111001000010100000000000;//SUB r[4],r[5] to r[7]
HD[2][70] <= 32'b10000000111000000000000000000000;//Output r[7]
HD[2][71] <= 32'b01110000000000000000000000000000;//Hlt
HD[2][72] <= 32'b00000000000000000000000000000000;
	 	 HD[2][128] <= 32'b01101100000000000000000000000000;//Nop
	 	 HD[2][129] <= 32'b01101000000000000000000000000000;//Loadi #0 to r[0]
	 	 HD[2][130] <= 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
	 	 HD[2][131] <= 32'b01101010110000000000000100000000;//Loadi #256 to r[22]
	 	 HD[2][132] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[2][133] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[2][134] <= 32'b01001100000000000000000000001010;//Branch on Zero #10
	 	 HD[2][135] <= 32'b10000111000101010000000000000000;//Loadr m[r[21]] to r[24]
	 	 HD[2][136] <= 32'b01011111001110000000000000000000;//SLT if r[24] < r[0], r[25] = 1 else r[25] = 0
	 	 HD[2][137] <= 32'b01011110111110011100000000000000;//SLT if r[25] < r[24], r[23] = 1 else r[23] = 0
	 	 HD[2][138] <= 32'b00100110111110011011100000000000;//OR r[25],r[23] to r[23]
	 	 HD[2][139] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[2][140] <= 32'b01001100000000000000000000000010;//Branch on Zero #2
	 	 HD[2][141] <= 32'b10000110111101010000000000000000;//Loadr m[r[21]] to r[23]
	 	 HD[2][142] <= 32'b10000010111000000000000000000000;//Output r[23]
	 	 HD[2][143] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[2][144] <= 32'b01010100000000000000000000000100;//Jump to #4
	 	 HD[2][145] <= 32'b01101010101000000000000000000000;//Loadi #0 to r[21]
	 	 HD[2][146] <= 32'b01101010110000000000000010010110;//Loadi #150 to r[22]
	 	 HD[2][147] <= 32'b01011110111101011011000000000000;//SLT if r[21] < r[22], r[23] = 1 else r[23] = 0
	 	 HD[2][148] <= 32'b01111100000101110000000000000000;//Pre Branch r[23]
	 	 HD[2][149] <= 32'b01001100000000000000000000001000;//Branch on Zero #8
	 	 HD[2][150] <= 32'b10000111000101010000000000000000;//Loadr m[r[21]] to r[24]
	 	 HD[2][151] <= 32'b01011111001000001100000000000000;//SLT if r[0] < r[24], r[25] = 1 else r[25] = 0
	 	 HD[2][152] <= 32'b01111100000110010000000000000000;//Pre Branch r[25]
	 	 HD[2][153] <= 32'b01001100000000000000000000000010;//Branch on Zero #2
	 	 HD[2][154] <= 32'b10010110111101010000000000000000;//LoadHD m[r[21]] to r[23]
	 	 HD[2][155] <= 32'b10000010111000000000000000000000;//Output r[23]
	 	 HD[2][156] <= 32'b00000110101101010000000000000001;//ADDi r[21], #1 to r[21]
	 	 HD[2][157] <= 32'b01010100000000000000000000010011;//Jump to #19
	 	 HD[2][158] <= 32'b01110000000000000000000000000000;//Hlt
		 HD[2][159] <= 32'b00000000000000000000000000000000;
		 HD[2][192] <= 32'b00000000000000000000000000000000;
			firstClock <= 1;
		end
	// Write
		if (flag_write_hd) begin
			HD[track][sector] <= data_write;
		end
	end


	// Continuous assignment implies read returns NEW data.
	// This is the natural behavior of the TriMatrix memory
	// blocks in Single Port mode.
	assign output_hard_drive = HD[track][sector];

endmodule
